
.subckt IVTRIX1_CV A C CN Y  BULKP BULKN AVDD AVSS
MN0 N1 A AVSS BULKN NCHDL
MN1 Y C N1 BULKN NCHDL
MP0 N2 A AVDD BULKP PCHDL
MP1 Y CN N2 BULKP PCHDL
.ends IVTRIX1_CV
