* CDAC8_CV 
.subckt CDAC8_CV  CP<11> CP<10> CP<9> CP<8> CP<7> CP<6> CP<5> CP<4> CP<3> CP<2> CP<1> CP<0> CTOP  AVSS
XC1  CP<10> CP<10> CP<10> CP<10> CP<10> CP<10> CTOP AVSS  CAP32C_CV
XC64a<0>  CP<8> CP<8> CP<8> CP<8> CP<8> CP<8> CTOP AVSS  CAP32C_CV
XC32a<0>  CP<6> CP<6> CP<6> CP<6> CP<6> CP<7> CTOP AVSS  CAP32C_CV
XCS       AVSS CP<0> CP<1> CP<2> CP<3>  AVSS CTOP AVSS  CAP32C_CV
XC128a<1>  CP<11> CP<11> CP<11> CP<11> CP<11> CP<11> CTOP AVSS  CAP32C_CV
XC128b<2>  CP<10> CP<10> CP<10> CP<10> CP<10> CP<10> CTOP AVSS  CAP32C_CV
X16ab       CP<5> CP<5> CP<5> CP<5> CP<4> AVSS CTOP AVSS  CAP32C_CV
XC64b<1>  CP<9> CP<9> CP<9> CP<9> CP<9> CP<9> CTOP AVSS  CAP32C_CV
XC0 CP<11> CP<11> CP<11> CP<11> CP<11> CP<11> CTOP AVSS  CAP32C_CV
.ENDS CDAC8_CV
