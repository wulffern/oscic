* SARBSSW_CV 
.SUBCKT SARBSSW_CV VI CK  VO1 VO2 AVDD AVSS
M1 VI GN VO1 AVSS NCHDLR
M2 VI GN VO1 AVSS NCHDLR
M3 VI GN VO1 AVSS NCHDLR
M4 VI GN VO1 AVSS NCHDLR
M5 VI TIE_L VO2 AVSS NCHDLR
M6 VI TIE_L VO2 AVSS NCHDLR
M7 VI TIE_L VO2 AVSS NCHDLR
M8 VI TIE_L VO2 AVSS NCHDLR

XA0a AVSS TAPCELL_CV
XA0 CK CKN AVDD AVSS IVX1_CV
XA3 CKN CSRC VI VS AVDD AVSS TGPD_CV
XA4 CKN CSRC GN GNG TIE_H AVDD AVSS SARBSSWCTRL_CV
XA1 TIE_H AVDD AVSS TIEH_CV
XA2 TIE_L AVDD AVSS TIEL_CV
XA5 AVSS TAPCELL_CV
XCAPB GNG VS CAPX1_CV M=9
XCAPC GNG VS CAPX1_CV M=9

.ENDS
