* SWX4_CV 
.subckt SWX4_CV A Y VREF AVSS
MN0 Y A AVSS AVSS NCHDL
MN1 AVSS A Y AVSS NCHDL
MN2 Y A AVSS AVSS NCHDL
MN3 AVSS A Y AVSS NCHDL
MP0 Y A VREF AVSS PCHDL
MP1 VREF A Y AVSS PCHDL
MP2 Y A VREF AVSS PCHDL
MP3 VREF A Y AVSS PCHDL
.ends SWX4_CV
