* CDAC6_CV 
.subckt CDAC6_CV CP<5>  CP<4> CP<3> CP<2> CP<1> CP<0> CTOP  AVSS
XC1       AVSS CP<0> CP<1> CP<2> CP<3> CP<4> CTOP AVSS  CAP32C_CV
XC0       AVSS CP<5> CP<5> CP<5> CP<5>  CP<5> CTOP AVSS  CAP32C_CV
.ENDS
