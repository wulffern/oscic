**********************************************************************
**        Copyright (c) 2017 Carsten Wulff Software, Norway
** *******************************************************************
** Created       : wulff at 2017-9-23
** *******************************************************************
**   This program is free software: you can redistribute it and/or modify
**   it under the terms of the GNU General Public License as published by
**   the Free Software Foundation, either version 3 of the License, or
**   (at your option) any later version.
**
**   This program is distributed in the hope that it will be useful,
**   but WITHOUT ANY WARRANTY; without even the implied warranty of
**   MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
**   GNU General Public License for more details.
**
**   You should have received a copy of the GNU General Public License
**   along with this program.  If not, see <http://www.gnu.org/licenses/>.
**********************************************************************

.subckt RGRN8X1_CV  D<7> D<6> D<5> D<4> D<3> D<2> D<1> D<0> CK RN Q<7> Q<6> Q<5> Q<4> Q<3> Q<2> Q<1> Q<0> AVDD AVSS
XA0 D<0> CK Q<0> RN NC0 BULKP BULKN AVDD AVSS DFRNQNX1_CV
XB1 D<1> CK Q<1> RN NC1 BULKP BULKN AVDD AVSS DFRNQNX1_CV
XC2 D<2> CK Q<2> RN NC2 BULKP BULKN AVDD AVSS DFRNQNX1_CV
XD3 D<3> CK Q<3> RN NC3 BULKP BULKN AVDD AVSS DFRNQNX1_CV
XE4 D<4> CK Q<4> RN NC4 BULKP BULKN AVDD AVSS DFRNQNX1_CV
XF5 D<5> CK Q<5> RN NC5 BULKP BULKN AVDD AVSS DFRNQNX1_CV
XG6 D<6> CK Q<6> RN NC6 BULKP BULKN AVDD AVSS DFRNQNX1_CV
XH7 D<7> CK Q<7> RN NC7 BULKP BULKN AVDD AVSS DFRNQNX1_CV
.ends


.SUBCKT SRGRN8X1_CV SI CK SO AVDD AVSS
+ D<0> RN SI
XI0 SI D<7> D<6> D<5> D<4> D<3> D<2> D<1> CK  RN  D<7> D<6> D<5> D<4> 
+ D<3> D<2> D<1> SO  AVDD AVSS  RGRN8X1_CV
.ENDS

