
.subckt DFRNQNX1_CV D CK RN Q QN BULKP BULKN AVDD AVSS
XA0 BULKP BULKN TAPCELL_CV
XA1 CK RN CKN BULKP BULKN AVDD AVSS NDX1_CV
XA2 CKN CKB BULKP BULKN AVDD AVSS IVX1_CV
XA3 D CKN CKB A0 BULKP BULKN AVDD AVSS IVTRIX1_CV
XA4 A1 CKB CKN A0 BULKP BULKN AVDD AVSS IVTRIX1_CV
XA5 A0 A1 BULKP BULKN AVDD AVSS IVX1_CV
XA6 A1 CKB CKN QN BULKP BULKN AVDD AVSS IVTRIX1_CV
XA7 Q CKN CKB RN QN BULKP BULKN AVDD AVSS NDTRIX1_CV
XA8 QN Q BULKP BULKN AVDD AVSS IVX1_CV
.ends
