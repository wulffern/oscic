* SWX2_CV 
.subckt SWX2_CV A Y VREF AVSS
MN0 Y A AVSS AVSS NCHDL
MN1 AVSS A Y AVSS NCHDL
MP0 Y A VREF AVSS PCHDL
MP1 VREF A Y AVSS PCHDL
.ends SWX2_CV
