* CDAC10L_CV 
.SUBCKT CDAC10L_CV  CP<15> CP<14> CP<13> CP<12> CP<11> CP<10> CP<9> CP<8> CP<7> CP<6> CP<5> CP<4> CP<3> CP<2> CP<1> CP<0> CTOP  AVSS

XDMA1       AVSS   AVSS   AVSS   AVSS   AVSS   AVSS   AVSS  AVSS  CDAC_C32_CV
XC1         CP<15> CP<15> CP<15> CP<15> CP<15> CP<15> CTOP  AVSS  CDAC_C32_CV
XCD2        CP<14> CP<14> CP<14> CP<14> CP<14> CP<14> CTOP  AVSS  CDAC_C32_CV
XCA512a<1>  CP<14> CP<14> CP<14> CP<14> CP<14> CP<14> CTOP  AVSS  CDAC_C32_CV
XD512b<1>   CP<15> CP<15> CP<15> CP<15> CP<15> CP<15> CTOP  AVSS  CDAC_C32_CV
XE256b<7>   CP<12> CP<12> CP<12> CP<12> CP<12> CP<12> CTOP  AVSS  CDAC_C32_CV
XF256a<7>   CP<13> CP<13> CP<13> CP<13> CP<13> CP<13> CTOP  AVSS  CDAC_C32_CV
XG128b<3>   CP<10> CP<10> CP<10> CP<10> CP<10> CP<10> CTOP  AVSS  CDAC_C32_CV
XH64a<0>    CP<8>  CP<8>  CP<8>  CP<8>  CP<8>  CP<8>  CTOP  AVSS  CDAC_C32_CV
XAA16a      CP<5>  CP<5>  CP<5>  CP<5>  CP<4>  AVSS   CTOP  AVSS  CDAC_C32_CV
XKS         AVSS   CP<0>  CP<1>  CP<2>  CP<3>  AVSS   CTOP  AVSS  CDAC_C32_CV
XL128a<1>   CP<11> CP<11> CP<11> CP<11> CP<11> CP<11> CTOP  AVSS  CDAC_C32_CV
XN256a<5>   CP<13> CP<13> CP<13> CP<13> CP<13> CP<13> CTOP  AVSS  CDAC_C32_CV
XM256b<5>   CP<12> CP<12> CP<12> CP<12> CP<12> CP<12> CTOP  AVSS  CDAC_C32_CV
XO512a<2>   CP<14> CP<14> CP<14> CP<14> CP<14> CP<14> CTOP  AVSS  CDAC_C32_CV
XP512b<2>   CP<15> CP<15> CP<15> CP<15> CP<15> CP<15> CTOP  AVSS  CDAC_C32_CV
XQ512a<3>   CP<14> CP<14> CP<14> CP<14> CP<14> CP<14> CTOP  AVSS  CDAC_C32_CV
XR512b<3>   CP<15> CP<15> CP<15> CP<15> CP<15> CP<15> CTOP  AVSS  CDAC_C32_CV
XS512a<4>   CP<14> CP<14> CP<14> CP<14> CP<14> CP<14> CTOP  AVSS  CDAC_C32_CV
XT512b<4>   CP<15> CP<15> CP<15> CP<15> CP<15> CP<15> CTOP  AVSS  CDAC_C32_CV
XU512a<5>   CP<14> CP<14> CP<14> CP<14> CP<14> CP<14> CTOP  AVSS  CDAC_C32_CV
XV512b<5>   CP<15> CP<15> CP<15> CP<15> CP<15> CP<15> CTOP  AVSS  CDAC_C32_CV
XX256b<2>   CP<12> CP<12> CP<12> CP<12> CP<12> CP<12> CTOP  AVSS  CDAC_C32_CV
XY256a<2>   CP<13> CP<13> CP<13> CP<13> CP<13> CP<13> CTOP  AVSS  CDAC_C32_CV
XZ128b<2>   CP<10> CP<10> CP<10> CP<10> CP<10> CP<10> CTOP  AVSS  CDAC_C32_CV
XIB32<0>    CP<7>  CP<7>  CP<7>  CP<7>  CP<7>  CP<6>  CTOP  AVSS  CDAC_C32_CV
XABC64b<1>  CP<9>  CP<9>  CP<9>  CP<9>  CP<9>  CP<9>  CTOP  AVSS  CDAC_C32_CV
XACC128a<0> CP<11> CP<11> CP<11> CP<11> CP<11> CP<11> CTOP  AVSS  CDAC_C32_CV
XADC256b<0> CP<12> CP<12> CP<12> CP<12> CP<12> CP<12> CTOP  AVSS  CDAC_C32_CV
XAEC256a<0> CP<13> CP<13> CP<13> CP<13> CP<13> CP<13> CTOP  AVSS  CDAC_C32_CV
XAGC512b<6> CP<15> CP<15> CP<15> CP<15> CP<15> CP<15> CTOP  AVSS  CDAC_C32_CV
XAFC512a<6> CP<14> CP<14> CP<14> CP<14> CP<14> CP<14> CTOP  AVSS  CDAC_C32_CV
XAHC512a<7> CP<14> CP<14> CP<14> CP<14> CP<14> CP<14> CTOP  AVSS  CDAC_C32_CV
XBA0        CP<15> CP<15> CP<15> CP<15> CP<15> CP<15> CTOP  AVSS  CDAC_C32_CV
XDMB2       AVSS   AVSS   AVSS   AVSS   AVSS   AVSS   AVSS  AVSS  CDAC_C32_CV
.ENDS CDAC10_CV
