* SARTWOS2OFFSET_CV 
.SUBCKT SARTWOS2OFFSET_CV CTR<5> CTR<4> CTR<3> CTR<2> CTR<1> CTR<0>
+ CTRL_N<4> CTRL_N<3> CTRL_N<2> CTRL_N<1> CTRL_N<0> CTRL_P<4> CTRL_P<3>
+ CTRL_P<2> CTRL_P<1> CTRL_P<0> AVDD AVSS

XXC3<0> CTR<0>  CTR5_N CTRL_N<0> AVDD AVSS NRX1_CV
XXC2<0> CTR5_N  CTR<0> CTRL_P<0> AVDD AVSS  ANX1_CV

XXC3<1> CTR<1>  CTR5_N CTRL_N<1> AVDD AVSS NRX1_CV
XXC1 CTR<5> CTR5_N AVDD AVSS   IVX1_CV
XXC2<1> CTR5_N  CTR<1> CTRL_P<1> AVDD AVSS ANX1_CV


XXC2<2> CTR5_N  CTR<2> CTRL_P<2> AVDD AVSS ANX1_CV

XXC3<2> CTR<2>  CTR5_N CTRL_N<2> AVDD AVSS NRX1_CV
XXC3<3> CTR<3>  CTR5_N CTRL_N<3> AVDD AVSS NRX1_CV
XXC2<3> CTR5_N  CTR<3> CTRL_P<3> AVDD AVSS ANX1_CV



XXC2<4> CTR5_N CTR<4> CTRL_P<4> AVDD AVSS  ANX1_CV
XXC3<4> CTR<4>  CTR5_N CTRL_N<4> AVDD AVSS NRX1_CV
XXC0 AVSS TAPCELL_CV


.ENDS
