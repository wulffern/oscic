**********************************************************************
**        Copyright (c) 2018 Carsten Wulff Software, Norway 
** *******************************************************************
** Created       : wulff at 2018-3-19
** *******************************************************************
**  The MIT License (MIT)
** 
**  Permission is hereby granted, free of charge, to any person obtaining a copy
**  of this software and associated documentation files (the "Software"), to deal
**  in the Software without restriction, including without limitation the rights
**  to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
**  copies of the Software, and to permit persons to whom the Software is
**  furnished to do so, subject to the following conditions:
** 
**  The above copyright notice and this permission notice shall be included in all
**  copies or substantial portions of the Software.
** 
**  THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
**  IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
**  FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
**  AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
**  LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
**  OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
**  SOFTWARE.
**  
**********************************************************************



.subckt TGPD_CV C A B BULKP BULKN AVDD AVSS
MN0 AVSS C CN BULKN NCHDL
MN1 B C AVSS BULKN NCHDL
MN2 A CN B BULKN NCHDL
MP0 AVDD C CN BULKP PCHDL
MP1_DMY B AVDD AVDD BULKP PCHDL
MP2 A C B BULKP PCHDL
.ends

.subckt SARBSSWCTRL_CV C GN GNG TIE_H  BULKP BULKN AVDD AVSS
MN0 N1 C AVSS BULKN NCHDL
MN1 GN TIE_H N1 BULKN NCHDL
MP0 GNG C GN BULKP PCHDL
MP1 AVDD GN GNG BULKP PCHDL
.ends

.SUBCKT SAREMX1_CV A  B EN ENO RST_N BULKP BULKN AVDD AVSS
MN0 N3 EN AM BULKN  NCHDL
MN1 N3 B AVSS BULKN  NCHDL
MN2 AVSS A N3 BULKN  NCHDL
MN3 ENO AM AVSS BULKN  NCHDL
MP0 AVDD RST_N AM BULKP PCHDL
MP1 N2 B ENO BULKP  PCHDL
MP2 N1 A N2 BULKP  PCHDL
MP3 AVDD AM N1 BULKP  PCHDL
.ENDS

.SUBCKT SARLTX1_CV A CHL RST_N EN LCK_N BULKP BULKN AVDD AVSS
MN0 N1 A AVSS BULKN  NCHDL
MN1 N3 LCK_N N1 BULKN  NCHDL
MN2 CHL EN N3 BULKN  NCHDL
MP0 NP2 RST_N AVDD BULKP PCHDL
MP1 NP1 RST_N NP2 BULKP PCHDL
MP2 CHL RST_N NP1 BULKP PCHDL
.ENDS

.SUBCKT SARCEX1_CV A B Y RST AVDD AVSS
MN0 N4 RST AVSS AVSS  NCHDL
MN1 AVSS RST N4 AVSS  NCHDL
MN2 N1 RST AVSS AVSS  NCHDL
MN3 Y RST N1 AVSS  NCHDL

MP0 N2 A Y AVSS PCHDL
MP1 AVDD A N2 AVSS PCHDL
MP2 N3 B AVDD AVSS PCHDL
MP3 Y B N3 AVSS PCHDL
.ENDS

.SUBCKT SARCMPHX1_CV CI CK CO VMR N1 N2 BULKP BULKN AVDD AVSS
MN0  N1 CK AVSS BULKN NCHDL
MN1  N2 CI N1   BULKN NCHDL
MN2  N1 CI N2   BULKN NCHDL
MN3  N2 CI N1   BULKN NCHDL
MN4  N1 CI N2   BULKN NCHDL
MN5  N2 CI N1   BULKN NCHDL
MN6  CO VMR N2   BULKN NCHDL

MP0  AVDD CK N1 BULKP PCHDL
MP1  N2 CK AVDD BULKP PCHDL
MP2  AVDD AVDD N2 BULKP PCHDL
MP3  CO CK AVDD BULKP PCHDL
MP4  AVDD VMR CO BULKP PCHDL
MP5  CO VMR AVDD BULKP PCHDL
MP6  AVDD VMR CO BULKP PCHDL
.ENDS SARCMPHX1_CV


.SUBCKT SARKICKHX1_CV CI CK CKN BULKP BULKN AVDD AVSS
MN0  N1 CKN AVSS BULKN NCHDL
MN1  N1 CI N1   BULKN NCHDL
MN2  N1 CI N1   BULKN NCHDL
MN3  N1 CI N1   BULKN NCHDL
MN4  N1 CI N1   BULKN NCHDL
MN5  N1 CI N1   BULKN NCHDL
MN6  AVDD CK N1   BULKN NCHDL

MP0  AVDD CKN N1 BULKP PCHDL
MP1_DMY AVDD AVDD AVDD BULKP PCHDL
MP2_DMY AVDD AVDD AVDD BULKP PCHDL
MP3_DMY AVDD AVDD AVDD BULKP PCHDL
MP4_DMY AVDD AVDD AVDD BULKP PCHDL
MP5_DMY AVDD AVDD AVDD BULKP PCHDL
MP6_DMY  AVDD AVDD AVDD BULKP PCHDL
.ENDS SARKICKHX1_CV

*-----------------------------------------------------------------------------
* SAR composite logic cells
*---------------------------------------------------------------------------


.SUBCKT SARBSSW_CV VI CK CKN TIE_L VO1 VO2 AVDD AVSS
M0 NCHDLRDMY
M1 VI GN VO1 AVSS NCHDLR
M2 VI GN VO1 AVSS NCHDLR
M3 VI GN VO1 AVSS NCHDLR
M4 VI GN VO1 AVSS NCHDLR
M5 VI TIE_L VO2 AVSS NCHDLR
M6 VI TIE_L VO2 AVSS NCHDLR
M7 VI TIE_L VO2 AVSS NCHDLR
M8 VI TIE_L VO2 AVSS NCHDLR
M9 NCHDLRDMY

XA0a DMY_CV
XA0 CK CKN AVSS AVSS AVDD AVSS IVX1_CV
XA3 CKN VI VS AVSS AVSS AVDD AVSS TGPD_CV
XA4 CKN GN GNG TIE_H AVSS AVSS AVDD AVSS SARBSSWCTRL_CV
XA1 TIE_H AVSS AVSS AVDD AVSS TIEH_CV
XA2 TIE_L AVSS AVSS AVDD AVSS TIEL_CV
XA5 AVSS TAPCELL_CV
XA6 DMY_CV
XCAPB GNG VS CAPX1_CV M=7
XCAPC GNG VS CAPX1_CV M=7

.ENDS

.SUBCKT SARCMPX1_CV CPI CNI CPO CNO CK_CMP CK_SAMPLE DONE AVDD AVSS
XA0a DMY_CV
XA0 AVSS TAPCELL_CV
XA1 CPI CK_B CK_N AVSS AVSS AVDD AVSS SARKICKHX1_CV
XA2 CPI CK_B CNO_I CPO_I N1 NC1 AVSS AVSS AVDD AVSS SARCMPHX1_CV
XA2a CPO_I CPO AVSS AVSS AVDD AVSS IVX4_CV
XA3a CNO_I CNO AVSS AVSS AVDD AVSS IVX4_CV
XA3 CNI CK_B CPO_I CNO_I N1 NC2 AVSS AVSS  AVDD AVSS SARCMPHX1_CV
XA4 CNI CK_B CK_N AVSS AVSS AVDD AVSS SARKICKHX1_CV
XA9 CK_N CK_B AVSS AVSS AVDD AVSS IVX1_CV
XA10 DONE_N CK_A CK_N AVSS AVSS AVDD AVSS NDX1_CV
XA11 CK_SAMPLE DONE DONE_N AVSS AVSS AVDD AVSS NRX1_CV
XA12 CK_CMP CK_A AVSS AVSS AVDD AVSS IVX1_CV
XA13 AVSS TAPCELL_CV
XA14 DMY_CV
.ENDS


.SUBCKT SARMRYX1_CV CMP_OP CMP_ON EN RST_N ENO CHL_OP CHL_ON AVDD AVSS
XA0 AVSS TAPCELL_CV
XA1 CMP_OP CMP_ON EN ENO RST_N AVSS AVSS AVDD AVSS SAREMX1_CV
XA2 ENO LCK_N AVSS AVSS AVDD AVSS IVX1_CV
XA4 CMP_OP CHL_OP RST_N EN LCK_N AVSS AVSS AVDD AVSS SARLTX1_CV
XA5 CMP_ON CHL_ON RST_N EN LCK_N AVSS AVSS AVDD AVSS SARLTX1_CV
.ENDS

.SUBCKT SARDIGX1_CV CMP_OP CMP_ON EN RST_N ENO CP0 CP1 CN0 CN1 VREF AVDD AVSS
XA1 CMP_OP CMP_ON EN RST_N ENO CHL_OP CHL_ON AVDD AVSS SARMRYX1_CV
XA2 CHL_ON CN1 VREF AVSS SWX2_CV
XA3 CN1 CP1 VREF AVSS SWX2_CV
XA4 CHL_OP CP0 VREF AVSS SWX2_CV
XA5 CP0 CN0 VREF AVSS SWX2_CV
XA6 AVSS TAPCELL_CV
.ENDS

.SUBCKT SARDIGEX2_CV CMP_OP CMP_ON EN RST_N ENO DONE CP0 CP1 CN0 CN1 CEIN CEO CKS VREF AVDD AVSS
XA0a DMY_CV
XA1 CMP_OP CMP_ON EN RST_N ENO CHL_OP CHL_ON  AVDD AVSS SARMRYX1_CV

XA2 CHL_ON CN1 VREF AVSS SWX2_CV
XA3 CN1 CP1 VREF AVSS SWX2_CV
XA4 CHL_OP CP0 VREF AVSS SWX2_CV
XA5 CP0 CN0 VREF AVSS SWX2_CV

XA6 CN0 CP1 CE CKS AVDD AVSS SARCEX1_CV
XA7 ENO ENO_N AVSS AVSS AVDD AVSS IVX1_CV
XA8 ENO_N DONE AVSS AVSS AVDD AVSS IVX1_CV
XA9 ENO_N CE CE1 AVSS AVSS AVDD AVSS NDX1_CV
XA10 CE1 CE1_N AVSS AVSS AVDD AVSS IVX1_CV
XA11 CE1_N CEIN CEO1 AVSS AVSS AVDD AVSS NRX1_CV
XA12 CEO1 CEO AVSS AVSS AVDD AVSS IVX1_CV
XA13 AVSS TAPCELL_CV
XA14 DMY_CV
.ENDS
