* STATECTRL_CV 
.SUBCKT STATECTRL_CV A ACT1_CMP_N ACT2_CMP_N AVDD AVSS B CK_CMP EN ENO RST_N
XMN1 NN3 EN AVSS AVSS  NCHDL
XMN2 NN4 B NN3 AVSS  NCHDL
XMN3 NN4 A NN3 AVSS  NCHDL
XMN4 AM EN NN4 AVSS  NCHDL

XMN5 NN1 AM AVSS AVSS  NCHDL
XMN6 NN2 AM NN1 AVSS  NCHDL
XMN7 ENO AM NN2 AVSS  NCHDL
XMN9 CK_CMP EN NN2 AVSS  NCHDL


XMP1 AM RST_N AVDD AVSS  PCHDL
XMP3 N2 B ENO AVSS  PCHDL
XMP2 N1 A N2 AVSS  PCHDL
XMP6 NP2 ACT1_CMP_N N1 AVSS  PCHDL
XMP7 N1 ACT2_CMP_N NP2 AVSS  PCHDL
XMP4 AVDD AM N1 AVSS  PCHDL

XMP8 CK_CMP ENO NP2 AVSS  PCHDL
XMP9 CK_CMP RST_N AVDD AVSS  PCHDL
.ENDS
