* SAROFFSETCAL_CV 
.SUBCKT SAROFFSETCAL_CV  CALOFFSET<5> CALOFFSET<4> CALOFFSET<3>  CALOFFSET<2> CALOFFSET<1> CALOFFSET<0> OFF_N OFF_P AVDD AVSS


XA1 OFF_P CTRL_P<4> CTRL_P<3> CTRL_P<2> CTRL_P<1> CTRL_P<0> AVSS SAROFFSETCAL_NCH_CV
XB1 OFF_N CTRL_N<4> CTRL_N<3> CTRL_N<2> CTRL_N<1> CTRL_N<0> AVSS SAROFFSETCAL_NCHR_CV

XI15  CALOFFSET<5> CALOFFSET<4> CALOFFSET<3> CALOFFSET<2>
+ CALOFFSET<1> CALOFFSET<0> CTRL_N<4> CTRL_N<3> CTRL_N<2> CTRL_N<1> CTRL_N<0>
+ CTRL_P<4> CTRL_P<3> CTRL_P<2> CTRL_P<1> CTRL_P<0>  AVDD AVSS SARTWOS2OFFSET_CV
.ENDS
