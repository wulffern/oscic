* CDAC9H_CV 
.SUBCKT CDAC9H_CV  CP<13> CP<12> CP<11> CP<10> CP<9> CP<8> CP<7> CP<6> CP<5> CP<4> CP<3> CP<2> CP<1> CP<0> CTOP  AVSS
XC1  CP<13> CP<13> CP<13> CP<13> CP<13> CP<13> CP<12> CTOP  AVSS  CAP64CH_CV
XC128b<3>  CP<10> CP<10> CP<10> CP<10> CP<10> CP<10> CP<11> CTOP  AVSS  CAP64CH_CV
XCS        AVSS   CP<0>  CP<1>  CP<2>  CP<3>  AVSS   AVSS   CTOP   AVSS  CAP64CH_CV
XC32a<0>   CP<6> CP<6> CP<6> CP<6> CP<6> CP<7> AVSS  CTOP AVSS  CAP64CH_CV
XC256b<5>  CP<12> CP<12> CP<12> CP<12> CP<12> CP<12> CP<13> CTOP  AVSS  CAP64CH_CV
XC256a<2>  CP<13> CP<13> CP<13> CP<13> CP<13> CP<13> CP<12> CTOP   AVSS  CAP64CH_CV
X16ab      CP<5> CP<5> CP<5> CP<5> CP<4> AVSS AVSS CTOP  AVSS  CAP64CH_CV
XC64a<0>   CP<8> CP<8> CP<8> CP<8> CP<8> CP<8> CP<9> CTOP AVSS  CAP64CH_CV
XC128a<0>  CP<11> CP<11> CP<11> CP<11> CP<11> CP<11> CP<10>  CTOP  AVSS  CAP64CH_CV
XC0  CP<12> CP<12> CP<12> CP<12> CP<12> CP<12> CP<13>  CTOP  AVSS  CAP64CH_CV
.ENDS CDAC9_CV
