* TAPCELLBLK_CV 
.SUBCKT TAPCELLBLK_CV BLK_N BLK_P
MN1 BLK_N BLK_N BLK_N BLK_N  NCHDL
MP1 BLK_P BLK_P BLK_P BLK_P  PCHDL
.ENDS
