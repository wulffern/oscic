*Testbench for inverter
*----------------------------------------------------------------------------
* OPTIONS
*----------------------------------------------------------------------------
.option method=gear gmin=1e-12 reltol=1e-6

*----------------------------------------------------------------------------
* PARAMETERS
*----------------------------------------------------------------------------

.param vdd=1.2
.param vcm = 0.4
.param input_freq = 1e5

.param risefall = 1n
.param pw = 100n
.param per = 200n

*----------------------------------------------------------------------------
* INCULDE
*----------------------------------------------------------------------------
.include ../../ciccreator/sim/aimspice_model.spi
.include ../../build/tb_stdlib.spice


*----------------------------------------------------------------------------
* DUT
*----------------------------------------------------------------------------
xinv A B AVDD AVSS IVX1_CV



*----------------------------------------------------------------------------
* FORCE
*----------------------------------------------------------------------------
VDD AVDD 0 dc vdd
VSS AVSS 0 dc 0

VA A 0 pulse(0 vdd 0 risefall risefall pw per) dc 0

*----------------------------------------------------------------------------
* ANALYSIS
*----------------------------------------------------------------------------
.tran 1n 10u

*----------------------------------------------------------------------------
* PLOTS AND EXTRACTS
*----------------------------------------------------------------------------
.plot v(A)
.plot v(B)



