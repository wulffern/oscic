* TGPD_CV 
.subckt TGPD_CV C CSRC A B AVDD AVSS
MN0 AVSS C CN AVSS NCHDL
MN1 B C AVSS AVSS NCHDL
MN2 A CN B AVSS NCHDL
MN3 CSRC CN B AVSS NCHDL

MP0 AVDD C CN AVSS PCHDL
MP1 CSRC CN AVDD AVSS PCHDL
MP2 A C B AVSS PCHDL
MP3 CSRC C B AVSS PCHDL
.ends
