* TAPCELLB_CV 
.SUBCKT TAPCELLB_CV AVSS AVDD
MN1 AVSS AVSS AVSS AVSS  NCHDL
MP1 AVDD AVDD AVDD AVDD  PCHDL
.ENDS
