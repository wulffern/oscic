* SARCMPRX1_CV 
.SUBCKT SARCMPRX1_CV CPI CNI CPIR CNIR CPO CNO CK_CMP CK_SAMPLE PWRUP EN DONE NC1 NC2  AVDD AVSS
XA0 AVSS TAPCELL_CV
XA9 CK_CMP CK_B AVDD AVSS IVX1_CV
XA10 CK_B CK_N AVDD AVSS IVX1_CV
XA1 CPI CK_B CK_N AVDD AVSS SARKICKHX1_CV
XA2 CPI CK_B CNO_I CPO_I N1 NC1 AVDD AVSS SARCMPHX1_CV
XA2b CPIR CK_B CNO_I CPO_I N1A NC1 AVDD AVSS SARCMPHX1_CV

XA2a CPO_I CPO AVDD AVSS IVX4_CV
XA3a CNO_I CNO AVDD AVSS IVX4_CV

XA3b CNIR CK_B CPO_I CNO_I N1A NC2 AVDD AVSS SARCMPHX1_CV
XA3 CNI CK_B CPO_I CNO_I N1 NC2 AVDD AVSS SARCMPHX1_CV
XA4 CNI CK_B CK_N AVDD AVSS SARKICKHX1_CV

XA11 PWRUP CK_SAMPLE RST  AVDD AVSS NDX1_CV
XA13 TIEH DONE RST NC3 NN1 AVDD AVSS  DFRNQNX1_CV
XA12 TIEH AVDD AVSS  TIEH_CV
XA14 NN1 RST EN AVDD AVSS  ANX1_CV
XA15 AVSS TAPCELL_CV
.ENDS
