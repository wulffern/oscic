**********************************************************************
**        Copyright (c) 2017 Carsten Wulff Software, Norway
** *******************************************************************
** Created       : wulff at 2017-5-14
** *******************************************************************
**   This program is free software: you can redistribute it and/or modify
**   it under the terms of the GNU General Public License as published by
**   the Free Software Foundation, either version 3 of the License, or
**   (at your option) any later version.
**
**   This program is distributed in the hope that it will be useful,
**   but WITHOUT ANY WARRANTY; without even the implied warranty of
**   MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
**   GNU General Public License for more details.
**
**   You should have received a copy of the GNU General Public License
**   along with this program.  If not, see <http://www.gnu.org/licenses/>.
**********************************************************************


.subckt TIEH_CV Y BULKP BULKN AVDD AVSS
MN0 A A AVSS BULKN NCHDL
MP0 Y A AVDD BULKP PCHDL
.ends

.subckt TIEL_CV Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS AVSS NCHDL
MP0 A A AVDD AVSS PCHDL
.ends TIEL_CV


.subckt IVX1_CV A Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS BULKN NCHDL
MP0 Y A AVDD BULKP PCHDL
.ends

.subckt IVX2_CV A Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS BULKN NCHDL
MN1 AVSS A Y BULKN NCHDL
MP0 Y A AVDD BULKP PCHDL
MP1 AVDD A Y BULKP PCHDL
.ends

.subckt IVX4_CV A Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS BULKN NCHDL
MN1 AVSS A Y BULKN NCHDL
MN2 Y A AVSS BULKN NCHDL
MN3 AVSS A Y BULKN NCHDL
MP0 Y A AVDD BULKP PCHDL
MP1 AVDD A Y BULKP PCHDL
MP2 Y A AVDD BULKP PCHDL
MP3 AVDD A Y BULKP PCHDL
.ends IVX4_CV

.subckt IVX8_CV A Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS BULKN NCHDL
MN1 AVSS A Y BULKN NCHDL
MN2 Y A AVSS BULKN NCHDL
MN3 AVSS A Y BULKN NCHDL
MN4 Y A AVSS BULKN NCHDL
MN5 AVSS A Y BULKN NCHDL
MN6 Y A AVSS BULKN NCHDL
MN7 AVSS A Y BULKN NCHDL
MP0 Y A AVDD BULKP PCHDL
MP1 AVDD A Y BULKP PCHDL
MP2 Y A AVDD BULKP PCHDL
MP3 AVDD A Y BULKP PCHDL
MP4 Y A AVDD BULKP PCHDL
MP5 AVDD A Y BULKP PCHDL
MP6 Y A AVDD BULKP PCHDL
MP7 AVDD A Y BULKP PCHDL
.ends IVX8_CV

.subckt BFX1_CV A Y BULKP BULKN AVDD AVSS
MN0 AVSS A B BULKN NCHDL
MN1 Y B AVSS BULKN NCHDL
MP0 AVDD A B BULKP PCHDL
MP1 Y B AVDD BULKP PCHDL
.ends BFX1_CV



*-----------------------------------------------------------------------------
* NAND/NOR
*-----------------------------------------------------------------------------

.subckt NRX1_CV A B Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS BULKN  NCHDL
MN1 AVSS B Y BULKN  NCHDL
MP0 N1 A AVDD BULKP PCHDL
MP1 Y B N1 BULKP PCHDL
.ends NRX1_CV

.subckt NDX1_CV A B Y BULKP BULKN AVDD AVSS
MN0 N1 A AVSS BULKN NCHDL
MN1 Y B N1 BULKN NCHDL
MP0 Y A AVDD BULKP PCHDL
MP1 AVDD B Y BULKP PCHDL
.ends NDX1_CV

.subckt ORX1_CV A B Y BULKP BULKN AVDD AVSS
XA1 A B YN BULKP BULKN AVDD AVSS  NRX1_CV
XA2 YN Y BULKP BULKN AVDD AVSS  IVX1_CV
.ends

.subckt ANX1_CV A B Y BULKP BULKN AVDD AVSS
XA1 A B YN BULKP BULKN AVDD AVSS NDX1_CV
XA2 YN Y BULKP BULKN AVDD AVSS IVX1_CV
.ends


.subckt IVTRIX1_CV A C CN Y  BULKP BULKN AVDD AVSS
MN0 N1 A AVSS BULKN NCHDL
MN1 Y C N1 BULKN NCHDL
MP0 N2 A AVDD BULKP PCHDL
MP1 Y CN N2 BULKP PCHDL
.ends IVTRIX1_CV

.subckt NDTRIX1_CV A C CN RN Y BULKP BULKN AVDD AVSS
MN2 N1 RN AVSS BULKN NCHDL
MN0 N2 A N1 BULKN NCHDL
MN1 Y C N2 BULKN NCHDL
MP2 AVDD RN N2 BULKP PCHDL
MP0 N2 A AVDD BULKP PCHDL
MP1 Y CN N2 BULKP PCHDL
.ends


.subckt DFRNQNX1_CV D CK RN Q QN BULKP BULKN AVDD AVSS
XA0 BULKP BULKN TAPCELL_CV
XA1 CK RN CKN BULKP BULKN AVDD AVSS NDX1_CV
XA2 CKN CKB BULKP BULKN AVDD AVSS IVX1_CV
XA3 D CKN CKB A0 BULKP BULKN AVDD AVSS IVTRIX1_CV
XA4 A1 CKB CKN A0 BULKP BULKN AVDD AVSS IVTRIX1_CV
XA5 A0 A1 BULKP BULKN AVDD AVSS IVX1_CV
XA6 A1 CKB CKN QN BULKP BULKN AVDD AVSS IVTRIX1_CV
XA7 Q CKN CKB RN QN BULKP BULKN AVDD AVSS NDTRIX1_CV
XA8 QN Q BULKP BULKN AVDD AVSS IVX1_CV
.ends


.SUBCKT SCX1_CV A Y BULKP BULKN  AVDD AVSS
XA2 N1 A AVSS BULKN  NCHDL
XA3 SCO A N1 BULKN  NCHDL
XA4a AVDD SCO N1 BULKN  NCHDL
XA4b AVDD SCO N1 BULKN  NCHDL
XA5 Y SCO AVSS BULKN  NCHDL

XB0 N2 A AVDD BULKP  PCHDL
XB1 SCO A N2 BULKP  PCHDL
XB3a N2 SCO AVSS BULKP  PCHDL
XB3b N2 SCO AVSS BULKP  PCHDL
XB4 Y SCO AVDD AVSS  PCHDL
.ends
