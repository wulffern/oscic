
.subckt IVX2_CV A Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS BULKN NCHDL
MN1 AVSS A Y BULKN NCHDL
MP0 Y A AVDD BULKP PCHDL
MP1 AVDD A Y BULKP PCHDL
.ends
