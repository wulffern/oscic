* SARCMPX1_CV 
.SUBCKT SARCMPX1_CV CPI CNI CPO CNO CK_CMP CK_SAMPLE DONE AVDD AVSS
XA0a DMY_CV
XA0 AVSS TAPCELL_CV
XA1 CPI CK_B CK_N AVSS AVSS AVDD AVSS SARKICKHX1_CV
XA2 CPI CK_B CNO_I CPO_I N1 NC1 AVSS AVSS AVDD AVSS SARCMPHX1_CV
XA2a CPO_I CPO AVSS AVSS AVDD AVSS IVX4_CV
XA3a CNO_I CNO AVSS AVSS AVDD AVSS IVX4_CV
XA3 CNI CK_B CPO_I CNO_I N1 NC2 AVSS AVSS  AVDD AVSS SARCMPHX1_CV
XA4 CNI CK_B CK_N AVSS AVSS AVDD AVSS SARKICKHX1_CV
XA9 CK_N CK_B AVSS AVSS AVDD AVSS IVX1_CV
XA10 DONE_N CK_A CK_N AVSS AVSS AVDD AVSS NDX1_CV
XA11 CK_SAMPLE DONE DONE_N AVSS AVSS AVDD AVSS NRX1_CV
XA12 CK_CMP CK_A AVSS AVSS AVDD AVSS IVX1_CV
XA13 AVSS TAPCELL_CV
XA14 DMY_CV
.ENDS
