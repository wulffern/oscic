* CAP64C_CV 
.subckt CAP64C_CV C1A C1B C2 C4 C8 C16 C32 CTOP AVSS
xr1 CTOP NCa
xr2 AVSS Ncb

xres1a C1A NC1 RM1
xres1b C1B NC2 RM1
xres2 C2 NC3 RM1
xres4 C4 NC4 RM1
xres8 C8 NC5 RM1
xres16 C16 NC6 RM1
xres32 C32 NC7 RM1
.ends
