* DLX1_CV 
.subckt DLX1_CV A Y AVDD AVSS
MN1 n1 A AVSS AVSS NCHDL
MN2a n2 A n1 AVSS NCHDL
MN2b n3a A n2 AVSS NCHDL
MN2c n3b A n3a AVSS NCHDL
MN2d n3 A n3b AVSS NCHDL
MN2e AN A n3 AVSS NCHDL
MN4 AVSS AVSS AN AVSS NCHDL
MN5 Y AN AVSS AVSS NCHDL

MP5 AVDD A AN AVSS PCHDL
MP1 np2 AN AVDD AVSS PCHDL
MP2a np3 AN np2 AVSS PCHDL
MP2b np4a AN np3 AVSS PCHDL
MP2c np4b AN np4a AVSS PCHDL
MP2d np4 AN np4b AVSS PCHDL
MP2e Y AN np4 AVSS PCHDL
MP4 AVDD AVDD Y AVSS PCHDL

.ends
