* SARNSCAPLOGIC_CV 
.SUBCKT SARNSCAPLOGIC_CV SARP SARN RESP RESN DONE_IN EN DONE_OUT AVDD AVSS

X0 AVSS TAPCELL_CV
X1a DONE_IN DN2 AVDD AVSS DLX1_CV
X1b DN2 DN3 AVDD AVSS DLX1_CV
X1c DN3 DN4 AVDD AVSS DLX1_CV
X1d DN4 DN5 AVDD AVSS DLX1_CV
X1e DN5 DLO AVDD AVSS DLX1_CV
X5 DONE_IN DLO DONE_OUT AVDD AVSS ANX1_CV
X5a DONE_IN EN SMPL AVDD AVSS ANX1_CV

X8 SARP SMPL RESP AVDD AVSS TGX2_CV
X9 SARN SMPL RESN AVDD AVSS TGX2_CV

X8a SARP TIEL RESN AVDD AVSS TGX2_CV
X9b SARN TIEL RESP AVDD AVSS TGX2_CV
X7 TIEL AVDD AVSS TIEL_CV

.ENDS
