
.subckt TIEL_CV Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS AVSS NCHDL
MP0 A A AVDD AVSS PCHDL
.ends TIEL_CV
