* SARDIGEX2_CV 
.SUBCKT SARDIGEX2_CV CMP_OP CMP_ON EN RST_N ENO ARST_N CP0 CP1 CN0 CN1 DO CK_CMP CK_SAMPLE VREF AVDD AVSS

XA0 AVSS TAPCELL_CV
XA1 CMP_OP CN0 CP1 AVDD AVSS CMP_ON CK_CMP EN ENO RST_N  STATECTRL_CV
XA2 ENO ENO_N AVDD AVSS  IVX1_CV

XA4 CMP_OP CHL_OP RST_N EN ENO_N AVDD AVSS SARLTX1_CV
XA5 CMP_ON CHL_ON RST_N EN ENO_N AVDD AVSS SARLTX1_CV

XA6 CHL_ON CN1 VREF AVSS SWX2_CV
XA7 CN1 CP1 VREF AVSS SWX2_CV

XA8 CHL_OP CP0 VREF AVSS SWX2_CV
XA9 CP0 CN0 VREF AVSS SWX2_CV

XA10 CP1 ENO ARST_N DINT net08 AVDD AVSS  DFRNQNX1_CV
XA11 DINT CK_SAMPLE ARST_N DO net015 AVDD AVSS  DFRNQNX1_CV
XA12 AVSS TAPCELL_CV
.ENDS
