* SARDIGEX2_CV 
.SUBCKT SARDIGEX2_CV CMP_OP CMP_ON EN RST_N ENO DONE CP0 CP1 CN0 CN1 CEIN CEO CKS VREF AVDD AVSS
XA0a DMY_CV
XA1 CMP_OP CMP_ON EN RST_N ENO CHL_OP CHL_ON  AVDD AVSS SARMRYX1_CV

XA2 CHL_ON CN1 VREF AVSS SWX2_CV
XA3 CN1 CP1 VREF AVSS SWX2_CV
XA4 CHL_OP CP0 VREF AVSS SWX2_CV
XA5 CP0 CN0 VREF AVSS SWX2_CV

XA6 CN0 CP1 CE CKS AVDD AVSS SARCEX1_CV
XA7 ENO ENO_N AVSS AVSS AVDD AVSS IVX1_CV
XA8 ENO_N DONE AVSS AVSS AVDD AVSS IVX1_CV
XA9 ENO_N CE CE1 AVSS AVSS AVDD AVSS NDX1_CV
XA10 CE1 CE1_N AVSS AVSS AVDD AVSS IVX1_CV
XA11 CE1_N CEIN CEO1 AVSS AVSS AVDD AVSS NRX1_CV
XA12 CEO1 CEO AVSS AVSS AVDD AVSS IVX1_CV
XA13 AVSS TAPCELL_CV
XA14 DMY_CV
.ENDS
