**********************************************************************
**        Copyright (c) 2017 Carsten Wulff Software, Norway 
** *******************************************************************
** Created       : wulff at 2017-6-24
** *******************************************************************
**   This program is free software: you can redistribute it and/or modify
**   it under the terms of the GNU General Public License as published by
**   the Free Software Foundation, either version 3 of the License, or
**   (at your option) any later version.
** 
**   This program is distributed in the hope that it will be useful,
**   but WITHOUT ANY WARRANTY; without even the implied warranty of
**   MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
**   GNU General Public License for more details.
** 
**   You should have received a copy of the GNU General Public License
**   along with this program.  If not, see <http://www.gnu.org/licenses/>.
**********************************************************************


.subckt SWX2_CV A Y VREF AVSS
MN0 Y A AVSS AVSS NCHDL
MN1 AVSS A Y AVSS NCHDL
MP0 Y A VREF AVSS PCHDL
MP1 VREF A Y AVSS PCHDL
.ends SWX2_CV

.subckt SWX4_CV A Y VREF AVSS
MN0 Y A AVSS AVSS NCHDL
MN1 AVSS A Y AVSS NCHDL
MN2 Y A AVSS AVSS NCHDL
MN3 AVSS A Y AVSS NCHDL
MP0 Y A VREF AVSS PCHDL
MP1 VREF A Y AVSS PCHDL
MP2 Y A VREF AVSS PCHDL
MP3 VREF A Y AVSS PCHDL
.ends SWX4_CV


.subckt TGX1_CV C A B BULKP BULKN AVDD AVSS
MN0 CN C AVSS BULKN NCHDL
MN1 A C B BULKN NCHDL
MP0 CN C AVDD BULKP PCHDL
MP1 A CN B BULKP PCHDL
.ends


.subckt TGX2_CV C A B BULKP BULKN AVDD AVSS
MN0 CN C AVSS BULKN NCHDL
MN1 A C B BULKN NCHDL
MN2 A C B BULKN NCHDL
MP0 CN C AVDD BULKP PCHDL
MP1 A CN B BULKP PCHDL
MP2 A CN B BULKP PCHDL
.ends




