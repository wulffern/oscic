* SARBSSWCTRL_CV 
.subckt SARBSSWCTRL_CV C GN GNG TIE_H  BULKP BULKN AVDD AVSS
MN0 N1 C AVSS BULKN NCHDL
MN1 GN TIE_H N1 BULKN NCHDL
MP0 GNG C GN BULKP PCHDL
MP1 AVDD GN GNG BULKP PCHDL
.ends
