* CDAC8L_CV 
.subckt CDAC8L_CV  CP<11> CP<10> CP<9> CP<8> CP<7> CP<6> CP<5> CP<4> CP<3> CP<2> CP<1> CP<0> CTOP  AVSS
XC1  CP<10> CP<10> CP<10> CP<10> CP<10> CP<10> CTOP AVSS  CDAC_C32_CV
XA64a<0>  CP<8> CP<8> CP<8> CP<8> CP<8> CP<8> CTOP AVSS  CDAC_C32_CV
XB32a<0>  CP<6> CP<6> CP<6> CP<6> CP<6> CP<7> CTOP AVSS  CDAC_C32_CV
XDS       AVSS CP<0> CP<1> CP<2> CP<3>  AVSS CTOP AVSS  CDAC_C32_CV

XE128a<1>  CP<11> CP<11> CP<11> CP<11> CP<11> CP<11> CTOP AVSS  CDAC_C32_CV
XF128b<2>  CP<10> CP<10> CP<10> CP<10> CP<10> CP<10> CTOP AVSS  CDAC_C32_CV

XG16ab       CP<5> CP<5> CP<5> CP<5> CP<4> AVSS CTOP AVSS  CDAC_C32_CV

XH64b<1>  CP<9> CP<9> CP<9> CP<9> CP<9> CP<9> CTOP AVSS  CDAC_C32_CV

XDMB10 CP<11> CP<11> CP<11> CP<11> CP<11> CP<11> CTOP AVSS  CDAC_C32_CV
.ENDS
