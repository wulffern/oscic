* SARMRYX1_CV 
.SUBCKT SARMRYX1_CV CMP_OP CMP_ON EN RST_N ENO CHL_OP CHL_ON AVDD AVSS
XA0 AVSS TAPCELL_CV
XA1 CMP_OP CMP_ON EN ENO RST_N AVSS AVSS AVDD AVSS SAREMX1_CV
XA2 ENO LCK_N AVSS AVSS AVDD AVSS IVX1_CV
XA4 CMP_OP CHL_OP RST_N EN LCK_N AVSS AVSS AVDD AVSS SARLTX1_CV
XA5 CMP_ON CHL_ON RST_N EN LCK_N AVSS AVSS AVDD AVSS SARLTX1_CV
.ENDS
