* SARBSSWCTRL_CV 
.subckt SARBSSWCTRL_CV C CSRC GN GNG TIE_H  AVDD AVSS
MN0 N1 C AVSS AVSS NCHDL
MN1 GN TIE_H N1 AVSS NCHDL
MP0 GNG CSRC GN AVSS PCHDL
MP1 AVDD GN GNG AVSS PCHDL
.ends
