* CDAC9L_CV 
.SUBCKT CDAC9L_CV  CP<13> CP<12> CP<11> CP<10> CP<9> CP<8> CP<7> CP<6> CP<5> CP<4> CP<3> CP<2> CP<1> CP<0> CTOP  AVSS
XDMA1       AVSS   AVSS   AVSS   AVSS   AVSS   AVSS   AVSS  AVSS  CDAC_C32_CV
XC1  CP<12> CP<12> CP<12> CP<12> CP<12> CP<12> CTOP AVSS  CDAC_C32_CV
XA256a<7>  CP<13> CP<13> CP<13> CP<13> CP<13> CP<13> CTOP AVSS  CDAC_C32_CV
XB128b<3>  CP<10> CP<10> CP<10> CP<10> CP<10> CP<10> CTOP AVSS  CDAC_C32_CV
XD64a<0>  CP<8> CP<8> CP<8> CP<8> CP<8> CP<8> CTOP AVSS  CDAC_C32_CV
XE32a<0>  CP<6> CP<6> CP<6> CP<6> CP<6> CP<7> CTOP AVSS  CDAC_C32_CV
XFS       AVSS CP<0> CP<1> CP<2> CP<3>  AVSS CTOP AVSS  CDAC_C32_CV
XH128a<1>  CP<11> CP<11> CP<11> CP<11> CP<11> CP<11> CTOP AVSS  CDAC_C32_CV
XI256b<5>  CP<12> CP<12> CP<12> CP<12> CP<12> CP<12> CTOP AVSS  CDAC_C32_CV
XJ256a<5>  CP<13> CP<13> CP<13> CP<13> CP<13> CP<13> CTOP AVSS  CDAC_C32_CV
XK256b<2>  CP<12> CP<12> CP<12> CP<12> CP<12> CP<12> CTOP AVSS  CDAC_C32_CV
XL256a<2>  CP<13> CP<13> CP<13> CP<13> CP<13> CP<13> CTOP AVSS  CDAC_C32_CV
XM128b<2>  CP<10> CP<10> CP<10> CP<10> CP<10> CP<10> CTOP AVSS  CDAC_C32_CV
XN16ab       CP<5> CP<5> CP<5> CP<5> CP<4> AVSS CTOP AVSS  CDAC_C32_CV
XO64b<1>  CP<9> CP<9> CP<9> CP<9> CP<9> CP<9> CTOP AVSS  CDAC_C32_CV
XP128a<0>  CP<11> CP<11> CP<11> CP<11> CP<11> CP<11> CTOP AVSS  CDAC_C32_CV
XQ256b<0>  CP<12> CP<12> CP<12> CP<12> CP<12> CP<12> CTOP AVSS  CDAC_C32_CV
XR0  CP<13> CP<13> CP<13> CP<13> CP<13> CP<13> CTOP AVSS  CDAC_C32_CV
XDMB1       AVSS   AVSS   AVSS   AVSS   AVSS   AVSS   AVSS  AVSS  CDAC_C32_CV
.ENDS
