* SARBSSW_CV 
.SUBCKT SARBSSW_CV VI CK CKN TIE_L VO1 VO2 AVDD AVSS
M0 NCHDLRDMY
M1 VI GN VO1 AVSS NCHDLR
M2 VI GN VO1 AVSS NCHDLR
M3 VI GN VO1 AVSS NCHDLR
M4 VI GN VO1 AVSS NCHDLR
M5 VI TIE_L VO2 AVSS NCHDLR
M6 VI TIE_L VO2 AVSS NCHDLR
M7 VI TIE_L VO2 AVSS NCHDLR
M8 VI TIE_L VO2 AVSS NCHDLR
M9 NCHDLRDMY

XA0a DMY_CV
XA0 CK CKN AVSS AVSS AVDD AVSS IVX1_CV
XA3 CKN VI VS AVSS AVSS AVDD AVSS TGPD_CV
XA4 CKN GN GNG TIE_H AVSS AVSS AVDD AVSS SARBSSWCTRL_CV
XA1 TIE_H AVSS AVSS AVDD AVSS TIEH_CV
XA2 TIE_L AVSS AVSS AVDD AVSS TIEL_CV
XA5 AVSS TAPCELL_CV
XA6 DMY_CV
XCAPB GNG VS CAPX1_CV M=7
XCAPC GNG VS CAPX1_CV M=7

.ENDS
