* RGRN8X1_CV 
.subckt RGRN8X1_CV  D<7> D<6> D<5> D<4> D<3> D<2> D<1> D<0> CK RN Q<7> Q<6> Q<5> Q<4> Q<3> Q<2> Q<1> Q<0> AVDD AVSS
XA0 D<0> CK Q<0> RN NC0 BULKP BULKN AVDD AVSS DFRNQNX1_CV
XB1 D<1> CK Q<1> RN NC1 BULKP BULKN AVDD AVSS DFRNQNX1_CV
XC2 D<2> CK Q<2> RN NC2 BULKP BULKN AVDD AVSS DFRNQNX1_CV
XD3 D<3> CK Q<3> RN NC3 BULKP BULKN AVDD AVSS DFRNQNX1_CV
XE4 D<4> CK Q<4> RN NC4 BULKP BULKN AVDD AVSS DFRNQNX1_CV
XF5 D<5> CK Q<5> RN NC5 BULKP BULKN AVDD AVSS DFRNQNX1_CV
XG6 D<6> CK Q<6> RN NC6 BULKP BULKN AVDD AVSS DFRNQNX1_CV
XH7 D<7> CK Q<7> RN NC7 BULKP BULKN AVDD AVSS DFRNQNX1_CV
.ends
