* SARDIGMX1_CV 
.SUBCKT SARDIGMX1_CV CMP_OP CMP_ON EN RST_N ENO ARST_N CP0 CN1  DO CK_CMP CK_SAMPLE VREF AVDD AVSS

XA0 AVSS TAPCELL_CV
XA1 CMP_OP CN0 CP1 AVDD AVSS CMP_ON CK_CMP EN ENO RST_N  STATECTRL_CV
XA2 ENO ENO_N AVDD AVSS  IVX1_CV
XA4 CMP_OP CHL_OP RST_N EN ENO_N AVDD AVSS SARLTX1_CV
XA5 CMP_ON CHL_ON RST_N EN ENO_N AVDD AVSS SARLTX1_CV

XA6 CHL_ON CN1 VREF AVSS SWX2_CV
XA8 CHL_OP CP0 VREF AVSS SWX2_CV
XA10 CP0 ENO ARST_N DO net08 AVDD AVSS  DFRNQNX1_CV

XA12 AVSS TAPCELL_CV
.ENDS
