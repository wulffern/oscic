* SAROFFSETCAL_NCH_CV 
.SUBCKT SAROFFSETCAL_NCH_CV OFF CTRL<4> CTRL<3> CTRL<2> CTRL<1> CTRL<0> AVSS

* XB0    OFF CTRL<0> OFF AVSS  NCHDL

* XB1<1> OFF CTRL<1> OFF AVSS  NCHDL
* XB1<0> OFF CTRL<1> OFF AVSS  NCHDL
* XB2<3> OFF CTRL<2> OFF AVSS  NCHDL
* XB2<2> OFF CTRL<2> OFF AVSS  NCHDL
* XB2<1> OFF CTRL<2> OFF AVSS  NCHDL
* XB2<0> OFF CTRL<2> OFF AVSS  NCHDL
* XB3<7> OFF CTRL<3> OFF AVSS  NCHDL
* XB3<6> OFF CTRL<3> OFF AVSS  NCHDL
* XB3<5> OFF CTRL<3> OFF AVSS  NCHDL
* XB3<4> OFF CTRL<3> OFF AVSS  NCHDL
* XB3<3> OFF CTRL<3> OFF AVSS  NCHDL
* XB3<2> OFF CTRL<3> OFF AVSS  NCHDL
* XB3<1> OFF CTRL<3> OFF AVSS  NCHDL
* XB3<0> OFF CTRL<3> OFF AVSS  NCHDL

* XB4<15> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<14> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<13> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<12> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<11> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<10> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<9> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<8> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<7> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<6> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<5> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<4> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<3> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<2> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<1> OFF CTRL<4> OFF AVSS  NCHDL
* XB4a OFF CTRL<4> OFF AVSS  NCHDL

XB0    NC6 CTRL<0> OFF AVSS  NCHDL

XB1<1> NC71 CTRL<1> OFF AVSS  NCHDL
XB1<0> NC72 CTRL<1> OFF AVSS  NCHDL
XB2<3> NC81 CTRL<2> OFF AVSS  NCHDL
XB2<2> NC82 CTRL<2> OFF AVSS  NCHDL
XB2<1> NC83 CTRL<2> OFF AVSS  NCHDL
XB2<0> NC84 CTRL<2> OFF AVSS  NCHDL
XB3<7> NC91 CTRL<3> OFF AVSS  NCHDL
XB3<6> NC92 CTRL<3> OFF AVSS  NCHDL
XB3<5> NC93 CTRL<3> OFF AVSS  NCHDL
XB3<4> NC94 CTRL<3> OFF AVSS  NCHDL
XB3<3> NC95 CTRL<3> OFF AVSS  NCHDL
XB3<2> NC96 CTRL<3> OFF AVSS  NCHDL
XB3<1> NC97 CTRL<3> OFF AVSS  NCHDL
XB3<0> NC98 CTRL<3> OFF AVSS  NCHDL

XB4<15> NC101 CTRL<4> OFF AVSS  NCHDL
XB4<14> NC102 CTRL<4> OFF AVSS  NCHDL
XB4<13> NC103 CTRL<4> OFF AVSS  NCHDL
XB4<12> NC104 CTRL<4> OFF AVSS  NCHDL
XB4<11> NC105 CTRL<4> OFF AVSS  NCHDL
XB4<10> NC106 CTRL<4> OFF AVSS  NCHDL
XB4<9> NC108 CTRL<4> OFF AVSS  NCHDL
XB4<8> NC109 CTRL<4> OFF AVSS  NCHDL
XB4<7> NC1010 CTRL<4> OFF AVSS  NCHDL
XB4<6> NC1011 CTRL<4> OFF AVSS  NCHDL
XB4<5> NC1012 CTRL<4> OFF AVSS  NCHDL
XB4<4> NC1013 CTRL<4> OFF AVSS  NCHDL
XB4<3> NC1014 CTRL<4> OFF AVSS  NCHDL
XB4<2> NC1015 CTRL<4> OFF AVSS  NCHDL
XB4<1> NC1016 CTRL<4> OFF AVSS  NCHDL
XB4a NC1017 CTRL<4> OFF AVSS  NCHDL

.ends
