* SARCMPHX1_CV 
.SUBCKT SARCMPHX1_CV CI CK CO VMR N1 N2 AVDD AVSS
MN0  N1 CK AVSS AVSS NCHDL
MN1  N2 CI N1   AVSS NCHDL
MN2  N1 CI N2   AVSS NCHDL
MN3  N2 CI N1   AVSS NCHDL
MN4  N1 CI N2   AVSS NCHDL
MN5  N2 CI N1   AVSS NCHDL
MN6  CO VMR N2   AVSS NCHDL

MP0  AVDD CK N1 AVSS PCHDL
MP1  N2 CK AVDD AVSS PCHDL
MP2  AVDD AVDD N2 AVSS PCHDL
MP3  CO CK AVDD AVSS PCHDL
MP4  AVDD VMR CO AVSS PCHDL
MP5  CO VMR AVDD AVSS PCHDL
MP6  AVDD VMR CO AVSS PCHDL
.ENDS SARCMPHX1_CV
