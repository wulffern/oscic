* CDAC11_CV 
.SUBCKT CDAC11_CV  CP<16> CP<17> CP<15> CP<14> CP<13> CP<12> CP<11> CP<10> CP<9> CP<8> CP<7> CP<6> CP<5> CP<4> CP<3> CP<2> CP<1> CP<0> CTOP  AVSS

XC1        CP<16> CP<16> CP<16> CP<16> CP<16> CP<16> CP<16> CTOP  AVSS  CAP64C_CV
XC1024<1>  CP<17> CP<17> CP<17> CP<17> CP<17> CP<17> CP<17> CTOP  AVSS  CAP64C_CV
XC1024<2>  CP<16> CP<16> CP<16> CP<16> CP<16> CP<16> CP<16> CTOP  AVSS  CAP64C_CV
XC1024<3>  CP<17> CP<17> CP<17> CP<17> CP<17> CP<17> CP<17> CTOP  AVSS  CAP64C_CV
XC512b<1>  CP<14> CP<14> CP<14> CP<14> CP<14> CP<14> CP<14> CTOP  AVSS  CAP64C_CV
XC512b<0>  CP<15> CP<15> CP<15> CP<15> CP<15> CP<15> CP<15> CTOP  AVSS  CAP64C_CV
XC256a<7>  CP<13> CP<13> CP<13> CP<13> CP<13> CP<13> CP<12> CTOP  AVSS  CAP64C_CV
XC128b<3>  CP<10> CP<10> CP<10> CP<10> CP<10> CP<10> CP<11> CTOP  AVSS  CAP64C_CV
XC32a<0>   CP<6> CP<6> CP<6> CP<6> CP<6> CP<7> AVSS  CTOP AVSS  CAP64C_CV
XCS        AVSS   CP<0>  CP<1>  CP<2>  CP<3>  AVSS   AVSS   CTOP   AVSS  CAP64C_CV
XC256b<5>  CP<12> CP<12> CP<12> CP<12> CP<12> CP<12> CP<13> CTOP  AVSS  CAP64C_CV
XC512a<2>  CP<14> CP<14> CP<14> CP<14> CP<14> CP<14> CP<14> CTOP  AVSS  CAP64C_CV
XC512b<3>  CP<15> CP<15> CP<15> CP<15> CP<15> CP<15> CP<15> CTOP  AVSS  CAP64C_CV
XC1024<4>  CP<16> CP<16> CP<16> CP<16> CP<16> CP<16> CP<16> CTOP  AVSS  CAP64C_CV
XC1024<5>  CP<17> CP<17> CP<17> CP<17> CP<17> CP<17> CP<17> CTOP  AVSS  CAP64C_CV
XC1024<6>  CP<16> CP<16> CP<16> CP<16> CP<16> CP<16> CP<16> CTOP  AVSS  CAP64C_CV
XC1024<7>  CP<17> CP<17> CP<17> CP<17> CP<17> CP<17> CP<17> CTOP  AVSS  CAP64C_CV
XC1024<8>  CP<16> CP<16> CP<16> CP<16> CP<16> CP<16> CP<16> CTOP  AVSS  CAP64C_CV
XC1024<9>  CP<17> CP<17> CP<17> CP<17> CP<17> CP<17> CP<17> CTOP  AVSS  CAP64C_CV
XC1024<10> CP<16> CP<16> CP<16> CP<16> CP<16> CP<16> CP<16> CTOP  AVSS  CAP64C_CV
XC1024<11> CP<17> CP<17> CP<17> CP<17> CP<17> CP<17> CP<17> CTOP  AVSS  CAP64C_CV
XC512a<5>  CP<14> CP<14> CP<14> CP<14> CP<14> CP<14> CP<14> CTOP   AVSS  CAP64C_CV
XC512b<5>  CP<15> CP<15> CP<15> CP<15> CP<15> CP<15> CP<15> CTOP   AVSS  CAP64C_CV
XC256a<2>  CP<13> CP<13> CP<13> CP<13> CP<13> CP<13> CP<12> CTOP   AVSS  CAP64C_CV
XC64a<0>   CP<8> CP<8> CP<8> CP<8> CP<8> CP<8> CP<9> CTOP AVSS  CAP64C_CV
X16ab      CP<5> CP<5> CP<5> CP<5> CP<4> AVSS AVSS CTOP  AVSS  CAP64C_CV
XC128a<0>  CP<11> CP<11> CP<11> CP<11> CP<11> CP<11> CP<10>  CTOP  AVSS  CAP64C_CV
XC256b<0>  CP<12> CP<12> CP<12> CP<12> CP<12> CP<12> CP<13>  CTOP  AVSS  CAP64C_CV
XC512a<7>  CP<14> CP<14> CP<14> CP<14> CP<14> CP<14> CP<14>  CTOP  AVSS  CAP64C_CV
XC512a<6>  CP<15> CP<15> CP<15> CP<15> CP<15> CP<15> CP<15>  CTOP  AVSS  CAP64C_CV
XC1024<12> CP<16> CP<16> CP<16> CP<16> CP<16> CP<16> CP<16> CTOP  AVSS  CAP64C_CV
XC1024<13> CP<17> CP<17> CP<17> CP<17> CP<17> CP<17> CP<17> CTOP  AVSS  CAP64C_CV
XC1024<14> CP<16> CP<16> CP<16> CP<16> CP<16> CP<16> CP<16> CTOP  AVSS  CAP64C_CV
XC0        CP<17> CP<17> CP<17> CP<17> CP<17> CP<17> CP<17> CTOP  AVSS  CAP64C_CV
.ENDS CDAC11_CV
