**********************************************************************
**        Copyright (c) 2018 Carsten Wulff Software, Norway 
** *******************************************************************
** Created       : wulff at 2018-3-19
** *******************************************************************
**  The MIT License (MIT)
** 
**  Permission is hereby granted, free of charge, to any person obtaining a copy
**  of this software and associated documentation files (the "Software"), to deal
**  in the Software without restriction, including without limitation the rights
**  to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
**  copies of the Software, and to permit persons to whom the Software is
**  furnished to do so, subject to the following conditions:
** 
**  The above copyright notice and this permission notice shall be included in all
**  copies or substantial portions of the Software.
** 
**  THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
**  IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
**  FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
**  AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
**  LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
**  OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
**  SOFTWARE.
**  
**********************************************************************
.subckt TGPD_CV C CSRC A B AVDD AVSS
MN0 AVSS C CN AVSS NCHDL
MN1 B C AVSS AVSS NCHDL
MN2 A CN B AVSS NCHDL
MN3 CSRC CN B AVSS NCHDL

MP0 AVDD C CN AVSS PCHDL
MP1 CSRC CN AVDD AVSS PCHDL
MP2 A C B AVSS PCHDL
MP3 CSRC C B AVSS PCHDL
.ends



.subckt IVTRIX1_CV A C CN Y AVDD AVSS
MN0 N1 A AVSS AVSS NCHDL
MN1 Y C N1 AVSS NCHDL
MP0 N2 A AVDD AVSS PCHDL
MP1 Y CN N2 AVSS PCHDL

.ends IVTRIX1_CV

.subckt NDTRIX1_CV A C CN RN Y AVDD AVSS
MN2 N1 RN AVSS AVSS NCHDL
MN0 N2 A N1 AVSS NCHDL
MN1 Y C N2 AVSS NCHDL
MP2 AVDD RN N2 AVSS PCHDL
MP0 N2 A AVDD AVSS PCHDL
MP1 Y CN N2 AVSS PCHDL
.ends

.subckt DFRNQNX1_CV D CK RN Q QN AVDD AVSS
XA1 CK RN CKN AVDD AVSS NDX1_CV
XA2 CKN CKB AVDD AVSS IVX1_CV
XA3 D CKN CKB A0 AVDD AVSS IVTRIX1_CV
XA4 A1 CKB CKN A0 AVDD AVSS IVTRIX1_CV
XA5 A0 A1 AVDD AVSS IVX1_CV
XA6 A1 CKB CKN QN AVDD AVSS IVTRIX1_CV
XA7 Q CKN CKB RN QN AVDD AVSS NDTRIX1_CV
XA8 QN Q AVDD AVSS IVX1_CV
.ends

.subckt SARBSSWCTRL_CV C CSRC GN GNG TIE_H  AVDD AVSS
MN0 N1 C AVSS AVSS NCHDL
MN1 GN TIE_H N1 AVSS NCHDL
MP0 GNG CSRC GN AVSS PCHDL
MP1 AVDD GN GNG AVSS PCHDL
.ends

.subckt SWX2_CV A Y VREF AVSS
MN0 Y A AVSS AVSS NCHDL
MN1 AVSS A Y AVSS NCHDL
MP0 Y A VREF AVSS PCHDL
MP1 VREF A Y AVSS PCHDL
.ends SWX2_CV

.SUBCKT TAPCELL_CV TAP
MN1 TAP TAP TAP TAP  NCHDL
MP1 TAP TAP TAP TAP  PCHDL
.ENDS

.SUBCKT TAPCELLBLK_CV BLK_N BLK_P
MN1 BLK_N BLK_N BLK_N BLK_N  NCHDL
MP1 BLK_P BLK_P BLK_P BLK_P  PCHDL
.ENDS

.SUBCKT TAPCELLB_CV AVSS AVDD
MN1 AVSS AVSS AVSS AVSS  NCHDL
MP1 AVDD AVDD AVDD AVDD  PCHDL
.ENDS

.subckt SWX4_CV A Y VREF AVSS
MN0 Y A AVSS AVSS NCHDL
MN1 AVSS A Y AVSS NCHDL
MN2 Y A AVSS AVSS NCHDL
MN3 AVSS A Y AVSS NCHDL
MP0 Y A VREF AVSS PCHDL
MP1 VREF A Y AVSS PCHDL
MP2 Y A VREF AVSS PCHDL
MP3 VREF A Y AVSS PCHDL
.ends IVX4_CV


.subckt TGX2_CV A C B AVDD AVSS
MN0 AVSS C CN AVSS NCHDL
MN5 A AVSS AVSS AVSS NCHDL
MN1 B C A AVSS NCHDL
MN2 A C B AVSS NCHDL
MN1b B C A AVSS NCHDL

MP0 AVDD C CN AVSS PCHDL
MP5 A AVDD AVDD AVSS PCHDL
MP1 B CN A AVSS PCHDL
MP2 A CN B AVSS PCHDL
MP1b B CN A AVSS PCHDL

.ends
.subckt DLX1_CV A Y AVDD AVSS
MN1 n1 A AVSS AVSS NCHDL
MN2a n2 A n1 AVSS NCHDL
MN2b n3a A n2 AVSS NCHDL
MN2c n3b A n3a AVSS NCHDL
MN2d n3 A n3b AVSS NCHDL
MN2e AN A n3 AVSS NCHDL
MN4 AVSS AVSS AN AVSS NCHDL
MN5 Y AN AVSS AVSS NCHDL

MP5 AVDD A AN AVSS PCHDL
MP1 np2 AN AVDD AVSS PCHDL
MP2a np3 AN np2 AVSS PCHDL
MP2b np4a AN np3 AVSS PCHDL
MP2c np4b AN np4a AVSS PCHDL
MP2d np4 AN np4b AVSS PCHDL
MP2e Y AN np4 AVSS PCHDL
MP4 AVDD AVDD Y AVSS PCHDL

.ends



*-----------------------------------------------------------------------------
* SAR unit logic cells
*---------------------------------------------------------------------------

.SUBCKT STATECTRL_CV A ACT1_CMP_N ACT2_CMP_N AVDD AVSS B CK_CMP EN ENO RST_N
XMN1 NN3 EN AVSS AVSS  NCHDL
XMN2 NN4 B NN3 AVSS  NCHDL
XMN3 NN4 A NN3 AVSS  NCHDL
XMN4 AM EN NN4 AVSS  NCHDL

XMN5 NN1 AM AVSS AVSS  NCHDL
XMN6 NN2 AM NN1 AVSS  NCHDL
XMN7 ENO AM NN2 AVSS  NCHDL
XMN9 CK_CMP EN NN2 AVSS  NCHDL


XMP1 AM RST_N AVDD AVSS  PCHDL
XMP3 N2 B ENO AVSS  PCHDL
XMP2 N1 A N2 AVSS  PCHDL
XMP6 NP2 ACT1_CMP_N N1 AVSS  PCHDL
XMP7 N1 ACT2_CMP_N NP2 AVSS  PCHDL
XMP4 AVDD AM N1 AVSS  PCHDL

XMP8 CK_CMP ENO NP2 AVSS  PCHDL
XMP9 CK_CMP RST_N AVDD AVSS  PCHDL
.ENDS


.SUBCKT SARLTX1_CV A CHL RST_N EN LCK_N AVDD AVSS
MN0 N1 A AVSS AVSS  NCHDL
MN1 N3 LCK_N N1 AVSS  NCHDL
MN2 CHL EN N3 AVSS  NCHDL
MP0 NP2 RST_N AVDD AVSS PCHDL
MP1 NP1 RST_N NP2 AVSS PCHDL
MP2 CHL RST_N NP1 AVSS PCHDL
.ENDS

.SUBCKT SARCMPHX1_CV CI CK CO VMR N1 N2 AVDD AVSS
MN0  N1 CK AVSS AVSS NCHDL
MN1  N2 CI N1   AVSS NCHDL
MN2  N1 CI N2   AVSS NCHDL
MN3  N2 CI N1   AVSS NCHDL
MN4  N1 CI N2   AVSS NCHDL
MN5  N2 CI N1   AVSS NCHDL
MN6  CO VMR N2   AVSS NCHDL

MP0  AVDD CK N1 AVSS PCHDL
MP1  N2 CK AVDD AVSS PCHDL
MP2  AVDD AVDD N2 AVSS PCHDL
MP3  CO CK AVDD AVSS PCHDL
MP4  AVDD VMR CO AVSS PCHDL
MP5  CO VMR AVDD AVSS PCHDL
MP6  AVDD VMR CO AVSS PCHDL
.ENDS SARCMPHX1_CV

.SUBCKT SARCMPHX0_CV CI CK CO VMR N1 N2 AVDD AVSS
MN0  N1 CK AVSS AVSS NCHDL
MN1  N2 CI N1   AVSS NCHDL
MN2  N1 CI N2   AVSS NCHDL
MN3  N2 CI N1   AVSS NCHDL
MN6  CO VMR N2   AVSS NCHDL

MP0  AVDD CK N1 AVSS PCHDL
MP1  N2 CK AVDD AVSS PCHDL

MP3  CO CK AVDD AVSS PCHDL
MP6  AVDD VMR CO AVSS PCHDL
.ENDS SARCMPHX1_CV

.SUBCKT SARKICKHX1_CV CI CK CKN AVDD AVSS
MN0  N1 CKN AVSS AVSS NCHDL
MN1  N1 CI N1   AVSS NCHDL
MN2  N1 CI N1   AVSS NCHDL
MN3  N1 CI N1   AVSS NCHDL
MN4  N1 CI N1   AVSS NCHDL
MN5  N1 CI N1   AVSS NCHDL
MN6  AVDD CK N1   AVSS NCHDL

MP0  AVDD CKN N1 AVSS PCHDL
MP1_DMY AVDD AVDD AVDD AVSS PCHDL
MP2_DMY AVDD AVDD AVDD AVSS PCHDL
MP3_DMY AVDD AVDD AVDD AVSS PCHDL
MP4_DMY AVDD AVDD AVDD AVSS PCHDL
MP5_DMY AVDD AVDD AVDD AVSS PCHDL
MP6  AVDD AVDD AVDD AVSS PCHDL
.ENDS SARKICKHX1_CV

*-----------------------------------------------------------------------------
* SAR composite logic cells
*---------------------------------------------------------------------------

.SUBCKT SARBSSW_CV VI CK  VO1 VO2 AVDD AVSS
M1 VI GN VO1 AVSS NCHDLR
M2 VI GN VO1 AVSS NCHDLR
M3 VI GN VO1 AVSS NCHDLR
M4 VI GN VO1 AVSS NCHDLR
M5 VI TIE_L VO2 AVSS NCHDLR
M6 VI TIE_L VO2 AVSS NCHDLR
M7 VI TIE_L VO2 AVSS NCHDLR
M8 VI TIE_L VO2 AVSS NCHDLR

XA0a AVSS TAPCELL_CV
XA0 CK CKN AVDD AVSS IVX1_CV
XA3 CKN CSRC VI VS AVDD AVSS TGPD_CV
XA4 CKN CSRC GN GNG TIE_H AVDD AVSS SARBSSWCTRL_CV
XA1 TIE_H AVDD AVSS TIEH_CV
XA2 TIE_L AVDD AVSS TIEL_CV
XA5 AVSS TAPCELL_CV
XCAPB GNG VS CAPX1_CV M=9
XCAPC GNG VS CAPX1_CV M=9

.ENDS

.SUBCKT SARCMPX0_CV CPI CNI CPO CNO CK_CMP CK_SAMPLE PWRUP EN DONE AVDD AVSS
XA0 AVSS TAPCELL_CV
XA9 CK_CMP CK_B AVDD AVSS IVX1_CV
XA10 CK_B CK_N AVDD AVSS IVX1_CV
XA2 CPI CK_B CNO_I CPO_I N1 NC1 AVDD AVSS SARCMPHX0_CV
XA2a CPO_I CPO AVDD AVSS IVX4_CV
XA3a CNO_I CNO AVDD AVSS IVX4_CV
XA3 CNI CK_B CPO_I CNO_I N1 NC2 AVDD AVSS SARCMPHX0_CV
XA11 PWRUP CK_SAMPLE RST  AVDD AVSS NDX1_CV
XA13 TIEH DONE RST NC3 NN1 AVDD AVSS  DFRNQNX1_CV
XA12 TIEH AVDD AVSS  TIEH_CV
XA14 NN1 RST EN AVDD AVSS  ANX1_CV
XA15 AVSS TAPCELL_CV
.ENDS

.SUBCKT SARCMPX1_CV CPI CNI CPO CNO CK_CMP CK_SAMPLE PWRUP EN DONE NC1 NC2 AVDD AVSS
XA0 AVSS TAPCELL_CV
XA9 CK_CMP CK_B AVDD AVSS IVX1_CV
XA10 CK_B CK_N AVDD AVSS IVX1_CV
XA1 CPI CK_B CK_N AVDD AVSS SARKICKHX1_CV
XA2 CPI CK_B CNO_I CPO_I N1 NC1 AVDD AVSS SARCMPHX1_CV

XA2a CPO_I CPO AVDD AVSS IVX4_CV
XA3a CNO_I CNO AVDD AVSS IVX4_CV

XA3 CNI CK_B CPO_I CNO_I N1 NC2 AVDD AVSS SARCMPHX1_CV
XA4 CNI CK_B CK_N AVDD AVSS SARKICKHX1_CV

XA11 PWRUP CK_SAMPLE RST  AVDD AVSS NDX1_CV
XA13 TIEH DONE RST NC3 NN1 AVDD AVSS  DFRNQNX1_CV
XA12 TIEH AVDD AVSS  TIEH_CV
XA14 NN1 RST EN AVDD AVSS  ANX1_CV
XA15 AVSS TAPCELL_CV
.ENDS

.SUBCKT SARCMPRX1_CV CPI CNI CPIR CNIR CPO CNO CK_CMP CK_SAMPLE PWRUP EN DONE NC1 NC2  AVDD AVSS
XA0 AVSS TAPCELL_CV
XA9 CK_CMP CK_B AVDD AVSS IVX1_CV
XA10 CK_B CK_N AVDD AVSS IVX1_CV
XA1 CPI CK_B CK_N AVDD AVSS SARKICKHX1_CV
XA2 CPI CK_B CNO_I CPO_I N1 NC1 AVDD AVSS SARCMPHX1_CV
XA2b CPIR CK_B CNO_I CPO_I N1A NC1 AVDD AVSS SARCMPHX1_CV

XA2a CPO_I CPO AVDD AVSS IVX4_CV
XA3a CNO_I CNO AVDD AVSS IVX4_CV

XA3b CNIR CK_B CPO_I CNO_I N1A NC2 AVDD AVSS SARCMPHX1_CV
XA3 CNI CK_B CPO_I CNO_I N1 NC2 AVDD AVSS SARCMPHX1_CV
XA4 CNI CK_B CK_N AVDD AVSS SARKICKHX1_CV

XA11 PWRUP CK_SAMPLE RST  AVDD AVSS NDX1_CV
XA13 TIEH DONE RST NC3 NN1 AVDD AVSS  DFRNQNX1_CV
XA12 TIEH AVDD AVSS  TIEH_CV
XA14 NN1 RST EN AVDD AVSS  ANX1_CV
XA15 AVSS TAPCELL_CV
.ENDS



.SUBCKT SARDIGEX2_CV CMP_OP CMP_ON EN RST_N ENO ARST_N CP0 CP1 CN0 CN1 DO CK_CMP CK_SAMPLE VREF AVDD AVSS

XA0 AVSS TAPCELL_CV
XA1 CMP_OP CN0 CP1 AVDD AVSS CMP_ON CK_CMP EN ENO RST_N  STATECTRL_CV
XA2 ENO ENO_N AVDD AVSS  IVX1_CV

XA4 CMP_OP CHL_OP RST_N EN ENO_N AVDD AVSS SARLTX1_CV
XA5 CMP_ON CHL_ON RST_N EN ENO_N AVDD AVSS SARLTX1_CV

XA6 CHL_ON CN1 VREF AVSS SWX2_CV
XA7 CN1 CP1 VREF AVSS SWX2_CV

XA8 CHL_OP CP0 VREF AVSS SWX2_CV
XA9 CP0 CN0 VREF AVSS SWX2_CV

XA10 CP1 ENO ARST_N DINT net08 AVDD AVSS  DFRNQNX1_CV
XA11 DINT CK_SAMPLE ARST_N DO net015 AVDD AVSS  DFRNQNX1_CV
XA12 AVSS TAPCELL_CV
.ENDS

.SUBCKT SARDIGMX1_CV CMP_OP CMP_ON EN RST_N ENO ARST_N CP0 CN1  DO CK_CMP CK_SAMPLE VREF AVDD AVSS

XA0 AVSS TAPCELL_CV
XA1 CMP_OP CN0 CP1 AVDD AVSS CMP_ON CK_CMP EN ENO RST_N  STATECTRL_CV
XA2 ENO ENO_N AVDD AVSS  IVX1_CV
XA4 CMP_OP CHL_OP RST_N EN ENO_N AVDD AVSS SARLTX1_CV
XA5 CMP_ON CHL_ON RST_N EN ENO_N AVDD AVSS SARLTX1_CV

XA6 CHL_ON CN1 VREF AVSS SWX2_CV
XA8 CHL_OP CP0 VREF AVSS SWX2_CV
XA10 CP0 ENO ARST_N DO net08 AVDD AVSS  DFRNQNX1_CV

XA12 AVSS TAPCELL_CV
.ENDS


.SUBCKT SARTWOS2OFFSET_CV CTR<5> CTR<4> CTR<3> CTR<2> CTR<1> CTR<0>
+ CTRL_N<4> CTRL_N<3> CTRL_N<2> CTRL_N<1> CTRL_N<0> CTRL_P<4> CTRL_P<3>
+ CTRL_P<2> CTRL_P<1> CTRL_P<0> AVDD AVSS

XXC3<0> CTR<0>  CTR5_N CTRL_N<0> AVDD AVSS NRX1_CV
XXC2<0> CTR5_N  CTR<0> CTRL_P<0> AVDD AVSS  ANX1_CV

XXC3<1> CTR<1>  CTR5_N CTRL_N<1> AVDD AVSS NRX1_CV
XXC1 CTR<5> CTR5_N AVDD AVSS   IVX1_CV
XXC2<1> CTR5_N  CTR<1> CTRL_P<1> AVDD AVSS ANX1_CV


XXC2<2> CTR5_N  CTR<2> CTRL_P<2> AVDD AVSS ANX1_CV

XXC3<2> CTR<2>  CTR5_N CTRL_N<2> AVDD AVSS NRX1_CV
XXC3<3> CTR<3>  CTR5_N CTRL_N<3> AVDD AVSS NRX1_CV
XXC2<3> CTR5_N  CTR<3> CTRL_P<3> AVDD AVSS ANX1_CV



XXC2<4> CTR5_N CTR<4> CTRL_P<4> AVDD AVSS  ANX1_CV
XXC3<4> CTR<4>  CTR5_N CTRL_N<4> AVDD AVSS NRX1_CV
XXC0 AVSS TAPCELL_CV


.ENDS

.SUBCKT SAROFFSETCAL_NCH_CV OFF CTRL<4> CTRL<3> CTRL<2> CTRL<1> CTRL<0> AVSS

* XB0    OFF CTRL<0> OFF AVSS  NCHDL

* XB1<1> OFF CTRL<1> OFF AVSS  NCHDL
* XB1<0> OFF CTRL<1> OFF AVSS  NCHDL
* XB2<3> OFF CTRL<2> OFF AVSS  NCHDL
* XB2<2> OFF CTRL<2> OFF AVSS  NCHDL
* XB2<1> OFF CTRL<2> OFF AVSS  NCHDL
* XB2<0> OFF CTRL<2> OFF AVSS  NCHDL
* XB3<7> OFF CTRL<3> OFF AVSS  NCHDL
* XB3<6> OFF CTRL<3> OFF AVSS  NCHDL
* XB3<5> OFF CTRL<3> OFF AVSS  NCHDL
* XB3<4> OFF CTRL<3> OFF AVSS  NCHDL
* XB3<3> OFF CTRL<3> OFF AVSS  NCHDL
* XB3<2> OFF CTRL<3> OFF AVSS  NCHDL
* XB3<1> OFF CTRL<3> OFF AVSS  NCHDL
* XB3<0> OFF CTRL<3> OFF AVSS  NCHDL

* XB4<15> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<14> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<13> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<12> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<11> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<10> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<9> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<8> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<7> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<6> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<5> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<4> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<3> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<2> OFF CTRL<4> OFF AVSS  NCHDL
* XB4<1> OFF CTRL<4> OFF AVSS  NCHDL
* XB4a OFF CTRL<4> OFF AVSS  NCHDL

XB0    NC6 CTRL<0> OFF AVSS  NCHDL

XB1<1> NC71 CTRL<1> OFF AVSS  NCHDL
XB1<0> NC72 CTRL<1> OFF AVSS  NCHDL
XB2<3> NC81 CTRL<2> OFF AVSS  NCHDL
XB2<2> NC82 CTRL<2> OFF AVSS  NCHDL
XB2<1> NC83 CTRL<2> OFF AVSS  NCHDL
XB2<0> NC84 CTRL<2> OFF AVSS  NCHDL
XB3<7> NC91 CTRL<3> OFF AVSS  NCHDL
XB3<6> NC92 CTRL<3> OFF AVSS  NCHDL
XB3<5> NC93 CTRL<3> OFF AVSS  NCHDL
XB3<4> NC94 CTRL<3> OFF AVSS  NCHDL
XB3<3> NC95 CTRL<3> OFF AVSS  NCHDL
XB3<2> NC96 CTRL<3> OFF AVSS  NCHDL
XB3<1> NC97 CTRL<3> OFF AVSS  NCHDL
XB3<0> NC98 CTRL<3> OFF AVSS  NCHDL

XB4<15> NC101 CTRL<4> OFF AVSS  NCHDL
XB4<14> NC102 CTRL<4> OFF AVSS  NCHDL
XB4<13> NC103 CTRL<4> OFF AVSS  NCHDL
XB4<12> NC104 CTRL<4> OFF AVSS  NCHDL
XB4<11> NC105 CTRL<4> OFF AVSS  NCHDL
XB4<10> NC106 CTRL<4> OFF AVSS  NCHDL
XB4<9> NC108 CTRL<4> OFF AVSS  NCHDL
XB4<8> NC109 CTRL<4> OFF AVSS  NCHDL
XB4<7> NC1010 CTRL<4> OFF AVSS  NCHDL
XB4<6> NC1011 CTRL<4> OFF AVSS  NCHDL
XB4<5> NC1012 CTRL<4> OFF AVSS  NCHDL
XB4<4> NC1013 CTRL<4> OFF AVSS  NCHDL
XB4<3> NC1014 CTRL<4> OFF AVSS  NCHDL
XB4<2> NC1015 CTRL<4> OFF AVSS  NCHDL
XB4<1> NC1016 CTRL<4> OFF AVSS  NCHDL
XB4a NC1017 CTRL<4> OFF AVSS  NCHDL

.ends


.SUBCKT SAROFFSETCAL_CV  CALOFFSET<5> CALOFFSET<4> CALOFFSET<3>  CALOFFSET<2> CALOFFSET<1> CALOFFSET<0> OFF_N OFF_P AVDD AVSS


XA1 OFF_P CTRL_P<4> CTRL_P<3> CTRL_P<2> CTRL_P<1> CTRL_P<0> AVSS SAROFFSETCAL_NCH_CV
XB1 OFF_N CTRL_N<4> CTRL_N<3> CTRL_N<2> CTRL_N<1> CTRL_N<0> AVSS SAROFFSETCAL_NCHR_CV

XI15  CALOFFSET<5> CALOFFSET<4> CALOFFSET<3> CALOFFSET<2>
+ CALOFFSET<1> CALOFFSET<0> CTRL_N<4> CTRL_N<3> CTRL_N<2> CTRL_N<1> CTRL_N<0>
+ CTRL_P<4> CTRL_P<3> CTRL_P<2> CTRL_P<1> CTRL_P<0>  AVDD AVSS SARTWOS2OFFSET_CV
.ENDS


.SUBCKT SARNSCAPLOGIC_CV SARP SARN RESP RESN DONE_IN EN DONE_OUT AVDD AVSS

X0 AVSS TAPCELL_CV
X1a DONE_IN DN2 AVDD AVSS DLX1_CV
X1b DN2 DN3 AVDD AVSS DLX1_CV
X1c DN3 DN4 AVDD AVSS DLX1_CV
X1d DN4 DN5 AVDD AVSS DLX1_CV
X1e DN5 DLO AVDD AVSS DLX1_CV
X5 DONE_IN DLO DONE_OUT AVDD AVSS ANX1_CV
X5a DONE_IN EN SMPL AVDD AVSS ANX1_CV

X8 SARP SMPL RESP AVDD AVSS TGX2_CV
X9 SARN SMPL RESN AVDD AVSS TGX2_CV

X8a SARP TIEL RESN AVDD AVSS TGX2_CV
X9b SARN TIEL RESP AVDD AVSS TGX2_CV
X7 TIEL AVDD AVSS TIEL_CV

.ENDS
