* IVTRIX1_CV 
.subckt IVTRIX1_CV A C CN Y AVDD AVSS
MN0 N1 A AVSS AVSS NCHDL
MN1 Y C N1 AVSS NCHDL
MP0 N2 A AVDD AVSS PCHDL
MP1 Y CN N2 AVSS PCHDL

.ends IVTRIX1_CV
