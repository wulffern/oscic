* CDAC_C32_CV 
.subckt CDAC_C32_CV C1A C1B C2 C4 C8 C16 CTOP AVSS

XA01  C16 CTOP AVSS CDAC_UNIT
XA02  C16 CTOP AVSS CDAC_UNIT
XA05  C8 CTOP AVSS CDAC_UNIT
XA03  C16 CTOP AVSS CDAC_UNIT
XA04  C16 CTOP AVSS CDAC_UNIT
XA06  C8 CTOP AVSS CDAC_UNIT

XA07  C4 CTOP AVSS CDAC_UNIT

XA08  C2 CTOP AVSS CDAC_UNIT

XA09  C1A CTOP AVSS CDAC_UNIT

XA10  C4 CTOP AVSS CDAC_UNIT

XA11  C8 CTOP AVSS CDAC_UNIT

XA13  C16 CTOP AVSS CDAC_UNIT
XA14  C16 CTOP AVSS CDAC_UNIT
XA12  C8 CTOP AVSS CDAC_UNIT
XA15  C16 CTOP AVSS CDAC_UNIT
XA16  C16 CTOP AVSS CDAC_UNIT

XA17  C16 CTOP AVSS CDAC_UNIT
XA18  C16 CTOP AVSS CDAC_UNIT
XA21  C8 CTOP AVSS CDAC_UNIT
XA19  C16 CTOP AVSS CDAC_UNIT
XA20  C16 CTOP AVSS CDAC_UNIT


XA22  C8 CTOP AVSS CDAC_UNIT

XA23  C4 CTOP AVSS CDAC_UNIT

XA24  C2 CTOP AVSS CDAC_UNIT

XA25  C1B CTOP AVSS CDAC_UNIT

XA26  C4 CTOP AVSS CDAC_UNIT

XA27  C8 CTOP AVSS CDAC_UNIT

XA29  C16 CTOP AVSS CDAC_UNIT
XA30  C16 CTOP AVSS CDAC_UNIT
XA28  C8 CTOP AVSS CDAC_UNIT
XA31  C16 CTOP AVSS CDAC_UNIT
XA32  C16 CTOP AVSS CDAC_UNIT
.ends
