* SARCEX1_CV 
.SUBCKT SARCEX1_CV A B Y RST AVDD AVSS
MN0 N4 RST AVSS AVSS  NCHDL
MN1 AVSS RST N4 AVSS  NCHDL
MN2 N1 RST AVSS AVSS  NCHDL
MN3 Y RST N1 AVSS  NCHDL

MP0 N2 A Y AVSS PCHDL
MP1 AVDD A N2 AVSS PCHDL
MP2 N3 B AVDD AVSS PCHDL
MP3 Y B N3 AVSS PCHDL
.ENDS
