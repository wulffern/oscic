* NDTRIX1_CV 
.subckt NDTRIX1_CV A C CN RN Y AVDD AVSS
MN2 N1 RN AVSS AVSS NCHDL
MN0 N2 A N1 AVSS NCHDL
MN1 Y C N2 AVSS NCHDL
MP2 AVDD RN N2 AVSS PCHDL
MP0 N2 A AVDD AVSS PCHDL
MP1 Y CN N2 AVSS PCHDL
.ends
