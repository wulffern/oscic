* TGX2_CV 
.subckt TGX2_CV A C B AVDD AVSS
MN0 AVSS C CN AVSS NCHDL
MN5 A AVSS AVSS AVSS NCHDL
MN1 B C A AVSS NCHDL
MN2 A C B AVSS NCHDL
MN1b B C A AVSS NCHDL

MP0 AVDD C CN AVSS PCHDL
MP5 A AVDD AVDD AVSS PCHDL
MP1 B CN A AVSS PCHDL
MP2 A CN B AVSS PCHDL
MP1b B CN A AVSS PCHDL

.ends
