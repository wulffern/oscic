* SARKICKHX1_CV 
.SUBCKT SARKICKHX1_CV CI CK CKN AVDD AVSS
MN0  N1 CKN AVSS AVSS NCHDL
MN1  N1 CI N1   AVSS NCHDL
MN2  N1 CI N1   AVSS NCHDL
MN3  N1 CI N1   AVSS NCHDL
MN4  N1 CI N1   AVSS NCHDL
MN5  N1 CI N1   AVSS NCHDL
MN6  AVDD CK N1   AVSS NCHDL

MP0  AVDD CKN N1 AVSS PCHDL
MP1_DMY AVDD AVDD AVDD AVSS PCHDL
MP2_DMY AVDD AVDD AVDD AVSS PCHDL
MP3_DMY AVDD AVDD AVDD AVSS PCHDL
MP4_DMY AVDD AVDD AVDD AVSS PCHDL
MP5_DMY AVDD AVDD AVDD AVSS PCHDL
MP6  AVDD AVDD AVDD AVSS PCHDL
.ENDS SARKICKHX1_CV
