* SARLTX1_CV 
.SUBCKT SARLTX1_CV A CHL RST_N EN LCK_N AVDD AVSS
MN0 N1 A AVSS AVSS  NCHDL
MN1 N3 LCK_N N1 AVSS  NCHDL
MN2 CHL EN N3 AVSS  NCHDL
MP0 NP2 RST_N AVDD AVSS PCHDL
MP1 NP1 RST_N NP2 AVSS PCHDL
MP2 CHL RST_N NP1 AVSS PCHDL
.ENDS
