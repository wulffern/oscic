* TAPCELL_CV 
.SUBCKT TAPCELL_CV TAP
MN1 TAP TAP TAP TAP  NCHDL
MP1 TAP TAP TAP TAP  PCHDL
.ENDS
