* SARDIGX1_CV 
.SUBCKT SARDIGX1_CV CMP_OP CMP_ON EN RST_N ENO CP0 CP1 CN0 CN1 VREF AVDD AVSS
XA1 CMP_OP CMP_ON EN RST_N ENO CHL_OP CHL_ON AVDD AVSS SARMRYX1_CV
XA2 CHL_ON CN1 VREF AVSS SWX2_CV
XA3 CN1 CP1 VREF AVSS SWX2_CV
XA4 CHL_OP CP0 VREF AVSS SWX2_CV
XA5 CP0 CN0 VREF AVSS SWX2_CV
XA6 AVSS TAPCELL_CV
.ENDS
