**********************************************************************
**        Copyright (c) 2017 Carsten Wulff Software, Norway 
** *******************************************************************
** Created       : wulff at 2017-6-11
** *******************************************************************
**   This program is free software: you can redistribute it and/or modify
**   it under the terms of the GNU General Public License as published by
**   the Free Software Foundation, either version 3 of the License, or
**   (at your option) any later version.
** 
**   This program is distributed in the hope that it will be useful,
**   but WITHOUT ANY WARRANTY; without even the implied warranty of
**   MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
**   GNU General Public License for more details.
** 
**   You should have received a copy of the GNU General Public License
**   along with this program.  If not, see <http://www.gnu.org/licenses/>.
**********************************************************************


.subckt CAPX A B D
XA  D A B  CAP M=10
.ends

.subckt CAPBW AIP AIN OTAIP OTAIN OTAOP OTAON AVSS
XB1 OTAON OTAIP AVSS CAPXT 
XB2 OTAON OTAIP AVSS CAPX yoffset=5 
XA1 OTAIP AIN AVSS CAPXT xoffset=5 
XA2 AIN OTAIN AVSS CAPX yoffset=5
XC1 OTAIN OTAOP AVSS CAPXT xoffset=5 
XC2 OTAIN OTAOP AVSS CAPX yoffset=5
.ends
