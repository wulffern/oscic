* CAPBW 
.subckt CAPBW AIP AIN OTAIP OTAIN OTAOP OTAON AVSS
XB1 OTAON OTAIP AVSS CAPXT 
XB2 OTAON OTAIP AVSS CAPX yoffset=5 
XA1 OTAIP AIN AVSS CAPXT xoffset=5 
XA2 AIN OTAIN AVSS CAPX yoffset=5
XC1 OTAIN OTAOP AVSS CAPXT xoffset=5 
XC2 OTAIN OTAOP AVSS CAPX yoffset=5
.ends
